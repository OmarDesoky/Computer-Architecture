LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY NewAddress IS
	PORT(PLA_ADDRESS : IN std_logic_vector(5 DOWNTO 0);		--ADDRESS FROM PLA
		BITOR_ADDRESS : IN std_logic_vector(5 DOWNTO 0);	--ADDRESS FROM BIT ORING
		 NEW_ADDRESS : OUT std_logic_vector(5 DOWNTO 0));	--OUTPUT NEW ADDRESS TO uAR

END ENTITY NewAddress;

ARCHITECTURE a_NewAddress OF NewAddress IS

BEGIN

	NEW_ADDRESS(0) <= PLA_ADDRESS(0) OR BITOR_ADDRESS(0);
	NEW_ADDRESS(1) <= PLA_ADDRESS(1) OR BITOR_ADDRESS(1);
	NEW_ADDRESS(2) <= PLA_ADDRESS(2) OR BITOR_ADDRESS(2);
	NEW_ADDRESS(3) <= PLA_ADDRESS(3) OR BITOR_ADDRESS(3);
	NEW_ADDRESS(4) <= PLA_ADDRESS(4) OR BITOR_ADDRESS(4);
	NEW_ADDRESS(5) <= PLA_ADDRESS(5) OR BITOR_ADDRESS(5);
	
END a_NewAddress;
